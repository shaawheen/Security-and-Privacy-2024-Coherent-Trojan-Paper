`ifndef DEVIL_REGISTER_FILE_VH
`define DEVIL_REGISTER_FILE_VH
`define DEVIL_REGISTER_FILE_CONTROL_EN_BIT_WIDTH 1
`define DEVIL_REGISTER_FILE_CONTROL_EN_BIT_MASK 1'h1
`define DEVIL_REGISTER_FILE_CONTROL_EN_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_CONTROL_TEST_BIT_WIDTH 4
`define DEVIL_REGISTER_FILE_CONTROL_TEST_BIT_MASK 4'hf
`define DEVIL_REGISTER_FILE_CONTROL_TEST_BIT_OFFSET 1
`define DEVIL_REGISTER_FILE_CONTROL_FUNC_BIT_WIDTH 4
`define DEVIL_REGISTER_FILE_CONTROL_FUNC_BIT_MASK 4'hf
`define DEVIL_REGISTER_FILE_CONTROL_FUNC_BIT_OFFSET 5
`define DEVIL_REGISTER_FILE_CONTROL_CRRESP_BIT_WIDTH 5
`define DEVIL_REGISTER_FILE_CONTROL_CRRESP_BIT_MASK 5'h1f
`define DEVIL_REGISTER_FILE_CONTROL_CRRESP_BIT_OFFSET 9
`define DEVIL_REGISTER_FILE_CONTROL_ACFLT_BIT_WIDTH 1
`define DEVIL_REGISTER_FILE_CONTROL_ACFLT_BIT_MASK 1'h1
`define DEVIL_REGISTER_FILE_CONTROL_ACFLT_BIT_OFFSET 14
`define DEVIL_REGISTER_FILE_CONTROL_ADDRFLT_BIT_WIDTH 1
`define DEVIL_REGISTER_FILE_CONTROL_ADDRFLT_BIT_MASK 1'h1
`define DEVIL_REGISTER_FILE_CONTROL_ADDRFLT_BIT_OFFSET 15
`define DEVIL_REGISTER_FILE_CONTROL_OSHEN_BIT_WIDTH 1
`define DEVIL_REGISTER_FILE_CONTROL_OSHEN_BIT_MASK 1'h1
`define DEVIL_REGISTER_FILE_CONTROL_OSHEN_BIT_OFFSET 16
`define DEVIL_REGISTER_FILE_CONTROL_CONEN_BIT_WIDTH 1
`define DEVIL_REGISTER_FILE_CONTROL_CONEN_BIT_MASK 1'h1
`define DEVIL_REGISTER_FILE_CONTROL_CONEN_BIT_OFFSET 17
`define DEVIL_REGISTER_FILE_CONTROL_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_CONTROL_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_CONTROL_BYTE_OFFSET 6'h00
`define DEVIL_REGISTER_FILE_STATUS_OSH_END_BIT_WIDTH 1
`define DEVIL_REGISTER_FILE_STATUS_OSH_END_BIT_MASK 1'h1
`define DEVIL_REGISTER_FILE_STATUS_OSH_END_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_STATUS_BUSY_BIT_WIDTH 1
`define DEVIL_REGISTER_FILE_STATUS_BUSY_BIT_MASK 1'h1
`define DEVIL_REGISTER_FILE_STATUS_BUSY_BIT_OFFSET 1
`define DEVIL_REGISTER_FILE_STATUS_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_STATUS_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_STATUS_BYTE_OFFSET 6'h04
`define DEVIL_REGISTER_FILE_DELAY_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_DELAY_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_DELAY_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_DELAY_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_DELAY_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_DELAY_BYTE_OFFSET 6'h08
`define DEVIL_REGISTER_FILE_ACSNOOP_TYPE_BIT_WIDTH 4
`define DEVIL_REGISTER_FILE_ACSNOOP_TYPE_BIT_MASK 4'hf
`define DEVIL_REGISTER_FILE_ACSNOOP_TYPE_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_ACSNOOP_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_ACSNOOP_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_ACSNOOP_BYTE_OFFSET 6'h0c
`define DEVIL_REGISTER_FILE_BASE_ADDR_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_BASE_ADDR_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_BASE_ADDR_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_BASE_ADDR_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_BASE_ADDR_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_BASE_ADDR_BYTE_OFFSET 6'h10
`define DEVIL_REGISTER_FILE_MEM_SIZE_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_MEM_SIZE_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_MEM_SIZE_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_MEM_SIZE_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_MEM_SIZE_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_MEM_SIZE_BYTE_OFFSET 6'h14
`define DEVIL_REGISTER_FILE_RDDATA_1_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_RDDATA_1_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_RDDATA_1_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_RDDATA_1_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_RDDATA_1_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_RDDATA_1_BYTE_OFFSET 6'h18
`define DEVIL_REGISTER_FILE_RDDATA_2_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_RDDATA_2_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_RDDATA_2_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_RDDATA_2_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_RDDATA_2_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_RDDATA_2_BYTE_OFFSET 6'h1c
`define DEVIL_REGISTER_FILE_RDDATA_3_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_RDDATA_3_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_RDDATA_3_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_RDDATA_3_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_RDDATA_3_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_RDDATA_3_BYTE_OFFSET 6'h20
`define DEVIL_REGISTER_FILE_RDDATA_4_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_RDDATA_4_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_RDDATA_4_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_RDDATA_4_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_RDDATA_4_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_RDDATA_4_BYTE_OFFSET 6'h24
`endif
