`ifndef DEVIL_REGISTER_FILE_VH
`define DEVIL_REGISTER_FILE_VH
`define DEVIL_REGISTER_FILE_CONTROL_EN_BIT_WIDTH 1
`define DEVIL_REGISTER_FILE_CONTROL_EN_BIT_MASK 1'h1
`define DEVIL_REGISTER_FILE_CONTROL_EN_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_CONTROL_TEST_BIT_WIDTH 4
`define DEVIL_REGISTER_FILE_CONTROL_TEST_BIT_MASK 4'hf
`define DEVIL_REGISTER_FILE_CONTROL_TEST_BIT_OFFSET 1
`define DEVIL_REGISTER_FILE_CONTROL_FUNC_BIT_WIDTH 4
`define DEVIL_REGISTER_FILE_CONTROL_FUNC_BIT_MASK 4'hf
`define DEVIL_REGISTER_FILE_CONTROL_FUNC_BIT_OFFSET 5
`define DEVIL_REGISTER_FILE_CONTROL_CRRESP_BIT_WIDTH 5
`define DEVIL_REGISTER_FILE_CONTROL_CRRESP_BIT_MASK 5'h1f
`define DEVIL_REGISTER_FILE_CONTROL_CRRESP_BIT_OFFSET 9
`define DEVIL_REGISTER_FILE_CONTROL_ACFLT_BIT_WIDTH 1
`define DEVIL_REGISTER_FILE_CONTROL_ACFLT_BIT_MASK 1'h1
`define DEVIL_REGISTER_FILE_CONTROL_ACFLT_BIT_OFFSET 14
`define DEVIL_REGISTER_FILE_CONTROL_ADDRFLT_BIT_WIDTH 1
`define DEVIL_REGISTER_FILE_CONTROL_ADDRFLT_BIT_MASK 1'h1
`define DEVIL_REGISTER_FILE_CONTROL_ADDRFLT_BIT_OFFSET 15
`define DEVIL_REGISTER_FILE_CONTROL_OSHEN_BIT_WIDTH 1
`define DEVIL_REGISTER_FILE_CONTROL_OSHEN_BIT_MASK 1'h1
`define DEVIL_REGISTER_FILE_CONTROL_OSHEN_BIT_OFFSET 16
`define DEVIL_REGISTER_FILE_CONTROL_CONEN_BIT_WIDTH 1
`define DEVIL_REGISTER_FILE_CONTROL_CONEN_BIT_MASK 1'h1
`define DEVIL_REGISTER_FILE_CONTROL_CONEN_BIT_OFFSET 17
`define DEVIL_REGISTER_FILE_CONTROL_ADLEN_BIT_WIDTH 1
`define DEVIL_REGISTER_FILE_CONTROL_ADLEN_BIT_MASK 1'h1
`define DEVIL_REGISTER_FILE_CONTROL_ADLEN_BIT_OFFSET 18
`define DEVIL_REGISTER_FILE_CONTROL_ADTEN_BIT_WIDTH 1
`define DEVIL_REGISTER_FILE_CONTROL_ADTEN_BIT_MASK 1'h1
`define DEVIL_REGISTER_FILE_CONTROL_ADTEN_BIT_OFFSET 19
`define DEVIL_REGISTER_FILE_CONTROL_PDTEN_BIT_WIDTH 1
`define DEVIL_REGISTER_FILE_CONTROL_PDTEN_BIT_MASK 1'h1
`define DEVIL_REGISTER_FILE_CONTROL_PDTEN_BIT_OFFSET 20
`define DEVIL_REGISTER_FILE_CONTROL_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_CONTROL_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_CONTROL_BYTE_OFFSET 8'h00
`define DEVIL_REGISTER_FILE_STATUS_OSH_END_BIT_WIDTH 1
`define DEVIL_REGISTER_FILE_STATUS_OSH_END_BIT_MASK 1'h1
`define DEVIL_REGISTER_FILE_STATUS_OSH_END_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_STATUS_BUSY_BIT_WIDTH 1
`define DEVIL_REGISTER_FILE_STATUS_BUSY_BIT_MASK 1'h1
`define DEVIL_REGISTER_FILE_STATUS_BUSY_BIT_OFFSET 1
`define DEVIL_REGISTER_FILE_STATUS_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_STATUS_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_STATUS_BYTE_OFFSET 8'h04
`define DEVIL_REGISTER_FILE_DELAY_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_DELAY_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_DELAY_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_DELAY_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_DELAY_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_DELAY_BYTE_OFFSET 8'h08
`define DEVIL_REGISTER_FILE_ACSNOOP_TYPE_BIT_WIDTH 4
`define DEVIL_REGISTER_FILE_ACSNOOP_TYPE_BIT_MASK 4'hf
`define DEVIL_REGISTER_FILE_ACSNOOP_TYPE_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_ACSNOOP_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_ACSNOOP_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_ACSNOOP_BYTE_OFFSET 8'h0c
`define DEVIL_REGISTER_FILE_BASE_ADDR_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_BASE_ADDR_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_BASE_ADDR_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_BASE_ADDR_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_BASE_ADDR_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_BASE_ADDR_BYTE_OFFSET 8'h10
`define DEVIL_REGISTER_FILE_MEM_SIZE_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_MEM_SIZE_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_MEM_SIZE_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_MEM_SIZE_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_MEM_SIZE_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_MEM_SIZE_BYTE_OFFSET 8'h14
`define DEVIL_REGISTER_FILE_ARSNOOP_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_ARSNOOP_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_ARSNOOP_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_ARSNOOP_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_ARSNOOP_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_ARSNOOP_BYTE_OFFSET 8'h18
`define DEVIL_REGISTER_FILE_L_ARADDR_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_L_ARADDR_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_L_ARADDR_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_L_ARADDR_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_L_ARADDR_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_L_ARADDR_BYTE_OFFSET 8'h1c
`define DEVIL_REGISTER_FILE_H_ARADDR_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_H_ARADDR_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_H_ARADDR_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_H_ARADDR_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_H_ARADDR_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_H_ARADDR_BYTE_OFFSET 8'h20
`define DEVIL_REGISTER_FILE_AWSNOOP_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_AWSNOOP_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_AWSNOOP_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_AWSNOOP_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_AWSNOOP_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_AWSNOOP_BYTE_OFFSET 8'h24
`define DEVIL_REGISTER_FILE_L_AWADDR_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_L_AWADDR_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_L_AWADDR_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_L_AWADDR_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_L_AWADDR_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_L_AWADDR_BYTE_OFFSET 8'h28
`define DEVIL_REGISTER_FILE_H_AWADDR_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_H_AWADDR_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_H_AWADDR_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_H_AWADDR_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_H_AWADDR_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_H_AWADDR_BYTE_OFFSET 8'h2c
`define DEVIL_REGISTER_FILE_RDATA_0_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_RDATA_0_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_RDATA_0_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_RDATA_0_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_RDATA_0_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_RDATA_0_BYTE_OFFSET 8'h40
`define DEVIL_REGISTER_FILE_WDATA_0_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_WDATA_0_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_WDATA_0_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_WDATA_0_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_WDATA_0_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_WDATA_0_BYTE_OFFSET 8'h40
`define DEVIL_REGISTER_FILE_RDATA_1_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_RDATA_1_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_RDATA_1_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_RDATA_1_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_RDATA_1_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_RDATA_1_BYTE_OFFSET 8'h44
`define DEVIL_REGISTER_FILE_WDATA_1_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_WDATA_1_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_WDATA_1_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_WDATA_1_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_WDATA_1_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_WDATA_1_BYTE_OFFSET 8'h44
`define DEVIL_REGISTER_FILE_RDATA_2_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_RDATA_2_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_RDATA_2_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_RDATA_2_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_RDATA_2_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_RDATA_2_BYTE_OFFSET 8'h48
`define DEVIL_REGISTER_FILE_WDATA_2_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_WDATA_2_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_WDATA_2_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_WDATA_2_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_WDATA_2_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_WDATA_2_BYTE_OFFSET 8'h48
`define DEVIL_REGISTER_FILE_RDATA_3_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_RDATA_3_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_RDATA_3_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_RDATA_3_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_RDATA_3_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_RDATA_3_BYTE_OFFSET 8'h4c
`define DEVIL_REGISTER_FILE_WDATA_3_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_WDATA_3_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_WDATA_3_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_WDATA_3_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_WDATA_3_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_WDATA_3_BYTE_OFFSET 8'h4c
`define DEVIL_REGISTER_FILE_RDATA_4_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_RDATA_4_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_RDATA_4_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_RDATA_4_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_RDATA_4_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_RDATA_4_BYTE_OFFSET 8'h50
`define DEVIL_REGISTER_FILE_WDATA_4_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_WDATA_4_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_WDATA_4_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_WDATA_4_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_WDATA_4_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_WDATA_4_BYTE_OFFSET 8'h50
`define DEVIL_REGISTER_FILE_RDATA_5_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_RDATA_5_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_RDATA_5_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_RDATA_5_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_RDATA_5_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_RDATA_5_BYTE_OFFSET 8'h54
`define DEVIL_REGISTER_FILE_WDATA_5_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_WDATA_5_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_WDATA_5_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_WDATA_5_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_WDATA_5_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_WDATA_5_BYTE_OFFSET 8'h54
`define DEVIL_REGISTER_FILE_RDATA_6_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_RDATA_6_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_RDATA_6_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_RDATA_6_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_RDATA_6_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_RDATA_6_BYTE_OFFSET 8'h58
`define DEVIL_REGISTER_FILE_WDATA_6_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_WDATA_6_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_WDATA_6_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_WDATA_6_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_WDATA_6_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_WDATA_6_BYTE_OFFSET 8'h58
`define DEVIL_REGISTER_FILE_RDATA_7_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_RDATA_7_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_RDATA_7_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_RDATA_7_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_RDATA_7_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_RDATA_7_BYTE_OFFSET 8'h5c
`define DEVIL_REGISTER_FILE_WDATA_7_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_WDATA_7_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_WDATA_7_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_WDATA_7_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_WDATA_7_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_WDATA_7_BYTE_OFFSET 8'h5c
`define DEVIL_REGISTER_FILE_RDATA_8_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_RDATA_8_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_RDATA_8_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_RDATA_8_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_RDATA_8_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_RDATA_8_BYTE_OFFSET 8'h60
`define DEVIL_REGISTER_FILE_WDATA_8_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_WDATA_8_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_WDATA_8_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_WDATA_8_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_WDATA_8_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_WDATA_8_BYTE_OFFSET 8'h60
`define DEVIL_REGISTER_FILE_RDATA_9_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_RDATA_9_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_RDATA_9_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_RDATA_9_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_RDATA_9_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_RDATA_9_BYTE_OFFSET 8'h64
`define DEVIL_REGISTER_FILE_WDATA_9_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_WDATA_9_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_WDATA_9_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_WDATA_9_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_WDATA_9_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_WDATA_9_BYTE_OFFSET 8'h64
`define DEVIL_REGISTER_FILE_RDATA_10_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_RDATA_10_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_RDATA_10_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_RDATA_10_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_RDATA_10_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_RDATA_10_BYTE_OFFSET 8'h68
`define DEVIL_REGISTER_FILE_WDATA_10_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_WDATA_10_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_WDATA_10_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_WDATA_10_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_WDATA_10_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_WDATA_10_BYTE_OFFSET 8'h68
`define DEVIL_REGISTER_FILE_RDATA_11_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_RDATA_11_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_RDATA_11_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_RDATA_11_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_RDATA_11_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_RDATA_11_BYTE_OFFSET 8'h6c
`define DEVIL_REGISTER_FILE_WDATA_11_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_WDATA_11_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_WDATA_11_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_WDATA_11_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_WDATA_11_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_WDATA_11_BYTE_OFFSET 8'h6c
`define DEVIL_REGISTER_FILE_RDATA_12_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_RDATA_12_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_RDATA_12_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_RDATA_12_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_RDATA_12_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_RDATA_12_BYTE_OFFSET 8'h70
`define DEVIL_REGISTER_FILE_WDATA_12_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_WDATA_12_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_WDATA_12_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_WDATA_12_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_WDATA_12_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_WDATA_12_BYTE_OFFSET 8'h70
`define DEVIL_REGISTER_FILE_RDATA_13_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_RDATA_13_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_RDATA_13_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_RDATA_13_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_RDATA_13_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_RDATA_13_BYTE_OFFSET 8'h74
`define DEVIL_REGISTER_FILE_WDATA_13_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_WDATA_13_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_WDATA_13_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_WDATA_13_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_WDATA_13_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_WDATA_13_BYTE_OFFSET 8'h74
`define DEVIL_REGISTER_FILE_RDATA_14_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_RDATA_14_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_RDATA_14_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_RDATA_14_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_RDATA_14_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_RDATA_14_BYTE_OFFSET 8'h78
`define DEVIL_REGISTER_FILE_WDATA_14_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_WDATA_14_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_WDATA_14_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_WDATA_14_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_WDATA_14_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_WDATA_14_BYTE_OFFSET 8'h78
`define DEVIL_REGISTER_FILE_RDATA_15_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_RDATA_15_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_RDATA_15_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_RDATA_15_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_RDATA_15_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_RDATA_15_BYTE_OFFSET 8'h7c
`define DEVIL_REGISTER_FILE_WDATA_15_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_WDATA_15_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_WDATA_15_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_WDATA_15_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_WDATA_15_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_WDATA_15_BYTE_OFFSET 8'h7c
`endif
