`ifndef DEVIL_REGISTER_FILE_VH
`define DEVIL_REGISTER_FILE_VH
`define DEVIL_REGISTER_FILE_CONTROL_EN_BIT_WIDTH 1
`define DEVIL_REGISTER_FILE_CONTROL_EN_BIT_MASK 1'h1
`define DEVIL_REGISTER_FILE_CONTROL_EN_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_CONTROL_TEST_BIT_WIDTH 4
`define DEVIL_REGISTER_FILE_CONTROL_TEST_BIT_MASK 4'hf
`define DEVIL_REGISTER_FILE_CONTROL_TEST_BIT_OFFSET 1
`define DEVIL_REGISTER_FILE_CONTROL_FUNC_BIT_WIDTH 4
`define DEVIL_REGISTER_FILE_CONTROL_FUNC_BIT_MASK 4'hf
`define DEVIL_REGISTER_FILE_CONTROL_FUNC_BIT_OFFSET 5
`define DEVIL_REGISTER_FILE_CONTROL_CRRESP_BIT_WIDTH 5
`define DEVIL_REGISTER_FILE_CONTROL_CRRESP_BIT_MASK 5'h1f
`define DEVIL_REGISTER_FILE_CONTROL_CRRESP_BIT_OFFSET 9
`define DEVIL_REGISTER_FILE_CONTROL_ACFLT_BIT_WIDTH 1
`define DEVIL_REGISTER_FILE_CONTROL_ACFLT_BIT_MASK 1'h1
`define DEVIL_REGISTER_FILE_CONTROL_ACFLT_BIT_OFFSET 14
`define DEVIL_REGISTER_FILE_CONTROL_ADDRFLT_BIT_WIDTH 1
`define DEVIL_REGISTER_FILE_CONTROL_ADDRFLT_BIT_MASK 1'h1
`define DEVIL_REGISTER_FILE_CONTROL_ADDRFLT_BIT_OFFSET 15
`define DEVIL_REGISTER_FILE_CONTROL_OSHEN_BIT_WIDTH 1
`define DEVIL_REGISTER_FILE_CONTROL_OSHEN_BIT_MASK 1'h1
`define DEVIL_REGISTER_FILE_CONTROL_OSHEN_BIT_OFFSET 16
`define DEVIL_REGISTER_FILE_CONTROL_CONEN_BIT_WIDTH 1
`define DEVIL_REGISTER_FILE_CONTROL_CONEN_BIT_MASK 1'h1
`define DEVIL_REGISTER_FILE_CONTROL_CONEN_BIT_OFFSET 17
`define DEVIL_REGISTER_FILE_CONTROL_ADLEN_BIT_WIDTH 1
`define DEVIL_REGISTER_FILE_CONTROL_ADLEN_BIT_MASK 1'h1
`define DEVIL_REGISTER_FILE_CONTROL_ADLEN_BIT_OFFSET 18
`define DEVIL_REGISTER_FILE_CONTROL_ADTEN_BIT_WIDTH 1
`define DEVIL_REGISTER_FILE_CONTROL_ADTEN_BIT_MASK 1'h1
`define DEVIL_REGISTER_FILE_CONTROL_ADTEN_BIT_OFFSET 19
`define DEVIL_REGISTER_FILE_CONTROL_PDTEN_BIT_WIDTH 1
`define DEVIL_REGISTER_FILE_CONTROL_PDTEN_BIT_MASK 1'h1
`define DEVIL_REGISTER_FILE_CONTROL_PDTEN_BIT_OFFSET 20
`define DEVIL_REGISTER_FILE_CONTROL_MONEN_BIT_WIDTH 1
`define DEVIL_REGISTER_FILE_CONTROL_MONEN_BIT_MASK 1'h1
`define DEVIL_REGISTER_FILE_CONTROL_MONEN_BIT_OFFSET 21
`define DEVIL_REGISTER_FILE_CONTROL_CMD_BIT_WIDTH 4
`define DEVIL_REGISTER_FILE_CONTROL_CMD_BIT_MASK 4'hf
`define DEVIL_REGISTER_FILE_CONTROL_CMD_BIT_OFFSET 22
`define DEVIL_REGISTER_FILE_CONTROL_BYTE_WIDTH 8
`define DEVIL_REGISTER_FILE_CONTROL_BYTE_SIZE 8
`define DEVIL_REGISTER_FILE_CONTROL_BYTE_OFFSET 9'h000
`define DEVIL_REGISTER_FILE_STATUS_OSH_END_BIT_WIDTH 1
`define DEVIL_REGISTER_FILE_STATUS_OSH_END_BIT_MASK 1'h1
`define DEVIL_REGISTER_FILE_STATUS_OSH_END_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_STATUS_BUSY_BIT_WIDTH 1
`define DEVIL_REGISTER_FILE_STATUS_BUSY_BIT_MASK 1'h1
`define DEVIL_REGISTER_FILE_STATUS_BUSY_BIT_OFFSET 1
`define DEVIL_REGISTER_FILE_STATUS_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_STATUS_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_STATUS_BYTE_OFFSET 9'h008
`define DEVIL_REGISTER_FILE_DELAY_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_DELAY_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_DELAY_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_DELAY_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_DELAY_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_DELAY_BYTE_OFFSET 9'h00c
`define DEVIL_REGISTER_FILE_ACSNOOP_TYPE_BIT_WIDTH 4
`define DEVIL_REGISTER_FILE_ACSNOOP_TYPE_BIT_MASK 4'hf
`define DEVIL_REGISTER_FILE_ACSNOOP_TYPE_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_ACSNOOP_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_ACSNOOP_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_ACSNOOP_BYTE_OFFSET 9'h010
`define DEVIL_REGISTER_FILE_BASE_ADDR_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_BASE_ADDR_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_BASE_ADDR_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_BASE_ADDR_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_BASE_ADDR_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_BASE_ADDR_BYTE_OFFSET 9'h014
`define DEVIL_REGISTER_FILE_MEM_SIZE_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_MEM_SIZE_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_MEM_SIZE_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_MEM_SIZE_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_MEM_SIZE_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_MEM_SIZE_BYTE_OFFSET 9'h018
`define DEVIL_REGISTER_FILE_ARSNOOP_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_ARSNOOP_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_ARSNOOP_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_ARSNOOP_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_ARSNOOP_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_ARSNOOP_BYTE_OFFSET 9'h01c
`define DEVIL_REGISTER_FILE_L_ARADDR_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_L_ARADDR_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_L_ARADDR_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_L_ARADDR_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_L_ARADDR_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_L_ARADDR_BYTE_OFFSET 9'h020
`define DEVIL_REGISTER_FILE_H_ARADDR_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_H_ARADDR_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_H_ARADDR_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_H_ARADDR_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_H_ARADDR_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_H_ARADDR_BYTE_OFFSET 9'h024
`define DEVIL_REGISTER_FILE_AWSNOOP_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_AWSNOOP_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_AWSNOOP_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_AWSNOOP_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_AWSNOOP_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_AWSNOOP_BYTE_OFFSET 9'h028
`define DEVIL_REGISTER_FILE_L_AWADDR_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_L_AWADDR_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_L_AWADDR_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_L_AWADDR_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_L_AWADDR_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_L_AWADDR_BYTE_OFFSET 9'h02c
`define DEVIL_REGISTER_FILE_H_AWADDR_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_H_AWADDR_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_H_AWADDR_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_H_AWADDR_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_H_AWADDR_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_H_AWADDR_BYTE_OFFSET 9'h030
`define DEVIL_REGISTER_FILE_RDATA_0_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_RDATA_0_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_RDATA_0_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_RDATA_0_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_RDATA_0_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_RDATA_0_BYTE_OFFSET 9'h040
`define DEVIL_REGISTER_FILE_WDATA_0_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_WDATA_0_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_WDATA_0_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_WDATA_0_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_WDATA_0_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_WDATA_0_BYTE_OFFSET 9'h040
`define DEVIL_REGISTER_FILE_RDATA_1_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_RDATA_1_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_RDATA_1_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_RDATA_1_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_RDATA_1_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_RDATA_1_BYTE_OFFSET 9'h044
`define DEVIL_REGISTER_FILE_WDATA_1_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_WDATA_1_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_WDATA_1_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_WDATA_1_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_WDATA_1_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_WDATA_1_BYTE_OFFSET 9'h044
`define DEVIL_REGISTER_FILE_RDATA_2_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_RDATA_2_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_RDATA_2_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_RDATA_2_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_RDATA_2_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_RDATA_2_BYTE_OFFSET 9'h048
`define DEVIL_REGISTER_FILE_WDATA_2_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_WDATA_2_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_WDATA_2_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_WDATA_2_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_WDATA_2_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_WDATA_2_BYTE_OFFSET 9'h048
`define DEVIL_REGISTER_FILE_RDATA_3_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_RDATA_3_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_RDATA_3_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_RDATA_3_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_RDATA_3_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_RDATA_3_BYTE_OFFSET 9'h04c
`define DEVIL_REGISTER_FILE_WDATA_3_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_WDATA_3_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_WDATA_3_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_WDATA_3_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_WDATA_3_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_WDATA_3_BYTE_OFFSET 9'h04c
`define DEVIL_REGISTER_FILE_RDATA_4_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_RDATA_4_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_RDATA_4_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_RDATA_4_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_RDATA_4_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_RDATA_4_BYTE_OFFSET 9'h050
`define DEVIL_REGISTER_FILE_WDATA_4_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_WDATA_4_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_WDATA_4_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_WDATA_4_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_WDATA_4_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_WDATA_4_BYTE_OFFSET 9'h050
`define DEVIL_REGISTER_FILE_RDATA_5_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_RDATA_5_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_RDATA_5_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_RDATA_5_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_RDATA_5_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_RDATA_5_BYTE_OFFSET 9'h054
`define DEVIL_REGISTER_FILE_WDATA_5_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_WDATA_5_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_WDATA_5_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_WDATA_5_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_WDATA_5_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_WDATA_5_BYTE_OFFSET 9'h054
`define DEVIL_REGISTER_FILE_RDATA_6_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_RDATA_6_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_RDATA_6_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_RDATA_6_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_RDATA_6_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_RDATA_6_BYTE_OFFSET 9'h058
`define DEVIL_REGISTER_FILE_WDATA_6_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_WDATA_6_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_WDATA_6_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_WDATA_6_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_WDATA_6_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_WDATA_6_BYTE_OFFSET 9'h058
`define DEVIL_REGISTER_FILE_RDATA_7_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_RDATA_7_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_RDATA_7_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_RDATA_7_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_RDATA_7_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_RDATA_7_BYTE_OFFSET 9'h05c
`define DEVIL_REGISTER_FILE_WDATA_7_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_WDATA_7_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_WDATA_7_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_WDATA_7_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_WDATA_7_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_WDATA_7_BYTE_OFFSET 9'h05c
`define DEVIL_REGISTER_FILE_RDATA_8_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_RDATA_8_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_RDATA_8_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_RDATA_8_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_RDATA_8_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_RDATA_8_BYTE_OFFSET 9'h060
`define DEVIL_REGISTER_FILE_WDATA_8_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_WDATA_8_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_WDATA_8_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_WDATA_8_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_WDATA_8_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_WDATA_8_BYTE_OFFSET 9'h060
`define DEVIL_REGISTER_FILE_RDATA_9_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_RDATA_9_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_RDATA_9_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_RDATA_9_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_RDATA_9_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_RDATA_9_BYTE_OFFSET 9'h064
`define DEVIL_REGISTER_FILE_WDATA_9_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_WDATA_9_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_WDATA_9_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_WDATA_9_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_WDATA_9_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_WDATA_9_BYTE_OFFSET 9'h064
`define DEVIL_REGISTER_FILE_RDATA_10_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_RDATA_10_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_RDATA_10_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_RDATA_10_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_RDATA_10_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_RDATA_10_BYTE_OFFSET 9'h068
`define DEVIL_REGISTER_FILE_WDATA_10_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_WDATA_10_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_WDATA_10_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_WDATA_10_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_WDATA_10_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_WDATA_10_BYTE_OFFSET 9'h068
`define DEVIL_REGISTER_FILE_RDATA_11_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_RDATA_11_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_RDATA_11_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_RDATA_11_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_RDATA_11_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_RDATA_11_BYTE_OFFSET 9'h06c
`define DEVIL_REGISTER_FILE_WDATA_11_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_WDATA_11_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_WDATA_11_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_WDATA_11_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_WDATA_11_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_WDATA_11_BYTE_OFFSET 9'h06c
`define DEVIL_REGISTER_FILE_RDATA_12_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_RDATA_12_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_RDATA_12_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_RDATA_12_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_RDATA_12_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_RDATA_12_BYTE_OFFSET 9'h070
`define DEVIL_REGISTER_FILE_WDATA_12_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_WDATA_12_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_WDATA_12_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_WDATA_12_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_WDATA_12_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_WDATA_12_BYTE_OFFSET 9'h070
`define DEVIL_REGISTER_FILE_RDATA_13_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_RDATA_13_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_RDATA_13_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_RDATA_13_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_RDATA_13_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_RDATA_13_BYTE_OFFSET 9'h074
`define DEVIL_REGISTER_FILE_WDATA_13_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_WDATA_13_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_WDATA_13_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_WDATA_13_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_WDATA_13_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_WDATA_13_BYTE_OFFSET 9'h074
`define DEVIL_REGISTER_FILE_RDATA_14_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_RDATA_14_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_RDATA_14_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_RDATA_14_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_RDATA_14_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_RDATA_14_BYTE_OFFSET 9'h078
`define DEVIL_REGISTER_FILE_WDATA_14_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_WDATA_14_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_WDATA_14_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_WDATA_14_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_WDATA_14_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_WDATA_14_BYTE_OFFSET 9'h078
`define DEVIL_REGISTER_FILE_RDATA_15_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_RDATA_15_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_RDATA_15_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_RDATA_15_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_RDATA_15_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_RDATA_15_BYTE_OFFSET 9'h07c
`define DEVIL_REGISTER_FILE_WDATA_15_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_WDATA_15_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_WDATA_15_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_WDATA_15_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_WDATA_15_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_WDATA_15_BYTE_OFFSET 9'h07c
`define DEVIL_REGISTER_FILE_PATTERN_0_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_PATTERN_0_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_PATTERN_0_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_PATTERN_0_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_PATTERN_0_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_PATTERN_0_BYTE_OFFSET 9'h080
`define DEVIL_REGISTER_FILE_PATTERN_1_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_PATTERN_1_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_PATTERN_1_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_PATTERN_1_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_PATTERN_1_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_PATTERN_1_BYTE_OFFSET 9'h084
`define DEVIL_REGISTER_FILE_PATTERN_2_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_PATTERN_2_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_PATTERN_2_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_PATTERN_2_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_PATTERN_2_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_PATTERN_2_BYTE_OFFSET 9'h088
`define DEVIL_REGISTER_FILE_PATTERN_3_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_PATTERN_3_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_PATTERN_3_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_PATTERN_3_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_PATTERN_3_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_PATTERN_3_BYTE_OFFSET 9'h08c
`define DEVIL_REGISTER_FILE_PATTERN_4_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_PATTERN_4_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_PATTERN_4_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_PATTERN_4_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_PATTERN_4_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_PATTERN_4_BYTE_OFFSET 9'h090
`define DEVIL_REGISTER_FILE_PATTERN_5_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_PATTERN_5_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_PATTERN_5_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_PATTERN_5_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_PATTERN_5_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_PATTERN_5_BYTE_OFFSET 9'h094
`define DEVIL_REGISTER_FILE_PATTERN_6_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_PATTERN_6_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_PATTERN_6_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_PATTERN_6_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_PATTERN_6_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_PATTERN_6_BYTE_OFFSET 9'h098
`define DEVIL_REGISTER_FILE_PATTERN_7_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_PATTERN_7_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_PATTERN_7_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_PATTERN_7_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_PATTERN_7_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_PATTERN_7_BYTE_OFFSET 9'h09c
`define DEVIL_REGISTER_FILE_PATTERN_8_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_PATTERN_8_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_PATTERN_8_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_PATTERN_8_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_PATTERN_8_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_PATTERN_8_BYTE_OFFSET 9'h0a0
`define DEVIL_REGISTER_FILE_PATTERN_9_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_PATTERN_9_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_PATTERN_9_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_PATTERN_9_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_PATTERN_9_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_PATTERN_9_BYTE_OFFSET 9'h0a4
`define DEVIL_REGISTER_FILE_PATTERN_10_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_PATTERN_10_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_PATTERN_10_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_PATTERN_10_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_PATTERN_10_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_PATTERN_10_BYTE_OFFSET 9'h0a8
`define DEVIL_REGISTER_FILE_PATTERN_11_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_PATTERN_11_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_PATTERN_11_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_PATTERN_11_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_PATTERN_11_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_PATTERN_11_BYTE_OFFSET 9'h0ac
`define DEVIL_REGISTER_FILE_PATTERN_12_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_PATTERN_12_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_PATTERN_12_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_PATTERN_12_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_PATTERN_12_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_PATTERN_12_BYTE_OFFSET 9'h0b0
`define DEVIL_REGISTER_FILE_PATTERN_13_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_PATTERN_13_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_PATTERN_13_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_PATTERN_13_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_PATTERN_13_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_PATTERN_13_BYTE_OFFSET 9'h0b4
`define DEVIL_REGISTER_FILE_PATTERN_14_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_PATTERN_14_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_PATTERN_14_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_PATTERN_14_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_PATTERN_14_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_PATTERN_14_BYTE_OFFSET 9'h0b8
`define DEVIL_REGISTER_FILE_PATTERN_15_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_PATTERN_15_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_PATTERN_15_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_PATTERN_15_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_PATTERN_15_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_PATTERN_15_BYTE_OFFSET 9'h0bc
`define DEVIL_REGISTER_FILE_PATTERN_SIZE_DATA_BIT_WIDTH 32
`define DEVIL_REGISTER_FILE_PATTERN_SIZE_DATA_BIT_MASK 32'hffffffff
`define DEVIL_REGISTER_FILE_PATTERN_SIZE_DATA_BIT_OFFSET 0
`define DEVIL_REGISTER_FILE_PATTERN_SIZE_BYTE_WIDTH 4
`define DEVIL_REGISTER_FILE_PATTERN_SIZE_BYTE_SIZE 4
`define DEVIL_REGISTER_FILE_PATTERN_SIZE_BYTE_OFFSET 9'h0c0
`endif
